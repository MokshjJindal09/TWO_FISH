`timescale 1ns / 1ps

module Mat_Multi(Key,S0,S1) ;
    input [127:0] Key;
    output [31:0] S0,S1;
    wire [7:0] S00,S01,S02,S03;
    wire [7:0] S10,S11,S12,S13;
    wire [7:0] A00,A01,A02,A03,A04,A05,A06,A07,A08,A09,A010,A011,A012,A013,A014,A015;
    wire [7:0] A10,A11,A12,A13,A14,A15,A16,A17,A18,A19,A110,A111,A112,A113,A114,A115;
    wire [7:0] A20,A21,A22,A23,A24,A25,A26,A27,A28,A29,A210,A211,A212,A213,A214,A215;
    wire [7:0] A30,A31,A32,A33,A34,A35,A36,A37,A38,A39,A310,A311,A312,A313,A314,A315;

    wire [7:0] m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,m15;
    
    assign {m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,m15} = Key;
    
    multi m000(8'h01,m0,9'b101001101,A00);
    multi m001(8'hA4,m1,9'b101001101,A01);
    multi m002(8'h55,m2,9'b101001101,A02);
    multi m003(8'h87,m3,9'b101001101,A03);
    multi m004(8'h5A,m4,9'b101001101,A04);
    multi m005(8'h58,m5,9'b101001101,A05);
    multi m006(8'hDB,m6,9'b101001101,A06);
    multi m007(8'h9E,m7,9'b101001101,A07);
    assign S00= A00^A01^A02^A03^A04^A05^A06^A07;


    multi m010(8'hA4,m0,9'b101001101,A10);
    multi m011(8'h56,m1,9'b101001101,A11);
    multi m012(8'h82,m2,9'b101001101,A12);
    multi m013(8'hF3,m3,9'b101001101,A13);
    multi m014(8'h1E,m4,9'b101001101,A14);
    multi m015(8'hC6,m5,9'b101001101,A15);
    multi m016(8'h68,m6,9'b101001101,A16);
    multi m017(8'hE5,m7,9'b101001101,A17);
    assign S01= A10^A11^A12^A13^A14^A15^A16^A17;


    multi m020(8'h02,m0,9'b101001101,A20);
    multi m021(8'hA1,m1,9'b101001101,A21);
    multi m022(8'hFC,m2,9'b101001101,A22);
    multi m023(8'hC1,m3,9'b101001101,A23);
    multi m024(8'h47,m4,9'b101001101,A24);
    multi m025(8'hAE,m5,9'b101001101,A25);
    multi m026(8'h3D,m6,9'b101001101,A26);
    multi m027(8'h19,m7,9'b101001101,A27);
    assign S02= A20^A21^A22^A23^A24^A25^A26^A27;


    multi m030(8'hA4,m0,9'b101001101,A30);
    multi m031(8'h55,m1,9'b101001101,A31);
    multi m032(8'h87,m2,9'b101001101,A32);
    multi m033(8'h5A,m3,9'b101001101,A33);
    multi m034(8'h58,m4,9'b101001101,A34);
    multi m035(8'hDB,m5,9'b101001101,A35);
    multi m036(8'h9E,m6,9'b101001101,A36);
    multi m037(8'h03,m7,9'b101001101,A37);
    assign S03= A30^A31^A32^A33^A34^A35^A36^A37;
    
    assign S1={S03,S02,S01,S00};
    
    
    
    
    
    multi m008(8'h01,m8,9'b101001101,A08);
    multi m009(8'hA4,m9,9'b101001101,A09);
    multi m0010(8'h55,m10,9'b101001101,A010);
    multi m0011(8'h87,m11,9'b101001101,A011);
    multi m0012(8'h5A,m12,9'b101001101,A012);
    multi m0013(8'h58,m13,9'b101001101,A013);
    multi m0014(8'hDB,m14,9'b101001101,A014);
    multi m0015(8'h9E,m15,9'b101001101,A015);
    assign S10= A08^A09^A010^A011^A012^A013^A014^A015;


    multi m018(8'hA4,m8,9'b101001101,A18);
    multi m019(8'h56,m9,9'b101001101,A19);
    multi m0110(8'h82,m10,9'b101001101,A110);
    multi m0111(8'hF3,m11,9'b101001101,A111);
    multi m0112(8'h1E,m12,9'b101001101,A112);
    multi m0113(8'hC6,m13,9'b101001101,A113);
    multi m0114(8'h68,m14,9'b101001101,A114);
    multi m0115(8'hE5,m15,9'b101001101,A115);
    assign S11= A18^A19^A110^A111^A112^A113^A114^A115;


    multi m028(8'h02,m8,9'b101001101,A28);
    multi m029(8'hA1,m9,9'b101001101,A29);
    multi m0210(8'hFC,m10,9'b101001101,A210);
    multi m0211(8'hC1,m11,9'b101001101,A211);
    multi m0212(8'h47,m12,9'b101001101,A212);
    multi m0213(8'hAE,m13,9'b101001101,A213);
    multi m0214(8'h3D,m14,9'b101001101,A214);
    multi m0215(8'h19,m15,9'b101001101,A215);
    assign S12= A28^A29^A210^A211^A212^A213^A214^A215;


    multi m038(8'hA4,m8,9'b101001101,A38);
    multi m039(8'h55,m9,9'b101001101,A39);
    multi m0310(8'h87,m10,9'b101001101,A310);
    multi m0311(8'h5A,m11,9'b101001101,A311);
    multi m0312(8'h58,m12,9'b101001101,A312);
    multi m0313(8'hDB,m13,9'b101001101,A313);
    multi m0314(8'h9E,m14,9'b101001101,A314);
    multi m0315(8'h03,m15,9'b101001101,A315);
    assign S13= A38^A39^A310^A311^A312^A313^A314^A315;
    
    assign S0={S13,S12,S11,S10};
endmodule